module judge3(
    input a,b,c,
    output out
);
    
    assign out = // 超过两个输入1
    
endmodule