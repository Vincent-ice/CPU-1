module timer(
	input clk,
    output [7:0] timer
);
    
    always @ (posedge clk) begin
    	...... 
    end
    
endmodule